module main

fn main() {
    
}