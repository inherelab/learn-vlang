module main

fn main() {
	println("hello vlang")
}
